//Design code
module w_or(
  input a,
  input b,
  output wor out);
  
  assign out = a ;
  assign out = b ;
  
endmodule
