//DESIGN CODE
module w_and(
  input a,
  input b,
  output wand out);
  
  assign out = a ;
  assign out = b ;
  
endmodule
