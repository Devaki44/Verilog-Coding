module diamond;
 initial begin
   $display("        1        ");
   $display("      2   2      ");
   $display("    3   3   3    ");
   $display("  4   4   4   4  ");
   $display("5   5   5   5   5");
   $display("  4   4   4   4  ");
   $display("    3   3   3    ");
   $display("      2   2      ");
   $display("        1        ");
 end
endmodule
